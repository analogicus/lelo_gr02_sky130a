** sch_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/BANDGAP/BANDGAP.sch
**.subckt BANDGAP VDD_1V8 I_PTAT V_CTAT PWRUP_1V8 VSS
*.ipin VDD_1V8
*.ipin VSS
*.opin I_PTAT
*.opin V_CTAT
*.ipin PWRUP_1V8
x1 VDD_1V8 PWRUP_1V8 V_B net2 V_CTAT VSS BANDGAP_OPAMP
x8 net1 PWRUP_1V8 VDD_1V8 VDD_1V8 JNWATR_PCH_12C1F2
x2 net2 V_B net1 VDD_1V8 JNWATR_PCH_4C1F2
x3 V_CTAT V_B net1 VDD_1V8 JNWATR_PCH_4C1F2
XQ1 VSS VSS net3 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=8 mult=8
XQ2 VSS VSS V_CTAT sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1 mult=1
x4 I_PTAT V_B net1 VDD_1V8 JNWATR_PCH_4C1F2
x5 net3 net2 VSS JNWTR_RPPO4
**.ends

* expanding   symbol:  BANDGAP_OPAMP/BANDGAP_OPAMP.sym # of pins=6
** sym_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/BANDGAP_OPAMP/BANDGAP_OPAMP.sym
** sch_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/BANDGAP_OPAMP/BANDGAP_OPAMP.sch
.subckt BANDGAP_OPAMP VDD_1V8 PWRUP_1V8 VOUT VIN_N VIN_P VSS
*.ipin VDD_1V8
*.ipin VSS
*.ipin PWRUP_1V8
*.ipin VIN_P
*.opin VOUT
*.ipin VIN_N
x8 SUPPLY PWRUP_1V8 VDD_1V8 VDD_1V8 JNWATR_PCH_12C1F2
R1 SUPPLY V_IB 100k m=1
x5<5> PMOS_GATE VIN_N TAIL VSS JNWATR_NCH_4C1F2
x5<4> PMOS_GATE VIN_N TAIL VSS JNWATR_NCH_4C1F2
x5<3> PMOS_GATE VIN_N TAIL VSS JNWATR_NCH_4C1F2
x5<2> PMOS_GATE VIN_N TAIL VSS JNWATR_NCH_4C1F2
x5<1> PMOS_GATE VIN_N TAIL VSS JNWATR_NCH_4C1F2
x5<0> PMOS_GATE VIN_N TAIL VSS JNWATR_NCH_4C1F2
x3<5> net1 VIN_P TAIL VSS JNWATR_NCH_4C1F2
x3<4> net1 VIN_P TAIL VSS JNWATR_NCH_4C1F2
x3<3> net1 VIN_P TAIL VSS JNWATR_NCH_4C1F2
x3<2> net1 VIN_P TAIL VSS JNWATR_NCH_4C1F2
x3<1> net1 VIN_P TAIL VSS JNWATR_NCH_4C1F2
x3<0> net1 VIN_P TAIL VSS JNWATR_NCH_4C1F2
x4 V_IB V_IB VSS VSS JNWATR_NCH_4C1F2
x6 TAIL V_IB VSS VSS JNWATR_NCH_4C1F2
x7 net1 PMOS_GATE SUPPLY VDD_1V8 JNWATR_PCH_4C1F2
x1 PMOS_GATE PMOS_GATE SUPPLY VDD_1V8 JNWATR_PCH_4C1F2
x2<2> VOUT net1 SUPPLY VDD_1V8 JNWATR_PCH_4C1F2
x2<1> VOUT net1 SUPPLY VDD_1V8 JNWATR_PCH_4C1F2
x2<0> VOUT net1 SUPPLY VDD_1V8 JNWATR_PCH_4C1F2
x3 VOUT V_IB VSS VSS JNWATR_NCH_4C1F2
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_PCH_12C1F2.sym # of pins=4
** sym_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_12C1F2.sym
** sch_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_12C1F2.sch
.subckt JNWATR_PCH_12C1F2 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.22 W=8.32 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_PCH_4C1F2.sym # of pins=4
** sym_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C1F2.sym
** sch_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C1F2.sch
.subckt JNWATR_PCH_4C1F2 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.22 W=3.2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RPPO4.sym # of pins=3
** sym_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO4.sym
** sch_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO4.sch
.subckt JNWTR_RPPO4 N P B
*.iopin P
*.iopin N
*.iopin B
XXA1 N P B JNWTR_RES4
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_NCH_4C1F2.sym # of pins=4
** sym_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_4C1F2.sym
** sch_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_4C1F2.sch
.subckt JNWATR_NCH_4C1F2 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.22 W=3.2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RES4.sym # of pins=3
** sym_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RES4.sym
** sch_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RES4.sch
.subckt JNWTR_RES4 N P B
*.iopin N
*.iopin P
*.iopin B
XR1_0 INT_0 N B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_1 INT_1 INT_0 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_2 INT_2 INT_1 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_3 P INT_2 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
.ends

.end
