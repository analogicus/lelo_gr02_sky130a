magic
tech sky130A
magscale 1 2
timestamp 1769081350
<< locali >>
rect 28516 21388 28834 21436
rect 28894 21388 28953 21436
rect 28516 21376 28953 21388
<< viali >>
rect 28834 21388 28894 21436
<< metal1 >>
rect 28834 21635 28894 21641
rect 28834 21442 28894 21575
rect 28822 21436 28906 21442
rect 28822 21388 28834 21436
rect 28894 21388 28906 21436
rect 28822 21382 28906 21388
<< via1 >>
rect 28834 21575 28894 21635
<< metal2 >>
rect 28834 21808 28894 21817
rect 28834 21635 28894 21752
rect 31864 21728 32132 21772
rect 29056 21723 31902 21728
rect 28828 21575 28834 21635
rect 28894 21575 28900 21635
rect 29052 21557 29061 21723
rect 29227 21557 31902 21723
rect 29056 21552 31902 21557
rect 32068 21552 32132 21728
rect 31864 21512 32132 21552
rect 31342 20788 31610 20826
rect 28516 20783 31386 20788
rect 28512 20617 28521 20783
rect 28687 20617 31386 20783
rect 28516 20612 31386 20617
rect 31552 20612 31610 20788
rect 31342 20566 31610 20612
rect 30705 13929 31095 13938
rect 30705 13530 31095 13539
rect 30205 13218 30595 13227
rect 30205 12819 30595 12828
rect 1104 11036 1113 11436
rect 1503 11036 1512 11436
rect 1634 10299 1643 10699
rect 2033 10299 2042 10699
<< via2 >>
rect 28834 21752 28894 21808
rect 29061 21557 29227 21723
rect 31902 21552 32068 21728
rect 28521 20617 28687 20783
rect 31386 20612 31552 20788
rect 30705 13539 31095 13929
rect 30205 12828 30595 13218
rect 1113 11036 1503 11436
rect 1643 10299 2033 10699
<< metal3 >>
rect 28832 21906 28896 21912
rect 28825 21842 28832 21895
rect 28896 21842 28916 21895
rect 28825 21808 28916 21842
rect 28825 21752 28834 21808
rect 28894 21752 28916 21808
rect 28825 21739 28916 21752
rect 31876 21733 32102 21764
rect 29056 21723 29232 21728
rect 29056 21557 29061 21723
rect 29227 21557 29232 21723
rect 29056 21310 29232 21557
rect 31876 21547 31897 21733
rect 32073 21547 32102 21733
rect 31876 21516 32102 21547
rect 28516 20783 28692 21022
rect 28516 20617 28521 20783
rect 28687 20617 28692 20783
rect 28516 20612 28692 20617
rect 31342 20793 31618 20840
rect 31342 20607 31381 20793
rect 31557 20607 31618 20793
rect 31342 20552 31618 20607
rect 30700 13929 31802 13934
rect 30700 13539 30705 13929
rect 31095 13539 31802 13929
rect 30700 13534 31802 13539
rect 32200 13534 32206 13934
rect 30200 13218 31323 13223
rect 30200 12828 30205 13218
rect 30595 12828 31323 13218
rect 30200 12823 31323 12828
rect 31721 12823 31727 13223
rect 1108 11436 1508 11441
rect -6 11036 0 11436
rect 398 11036 1113 11436
rect 1503 11036 1508 11436
rect 1108 11031 1508 11036
rect 1638 10699 2038 10704
rect 473 10299 479 10699
rect 877 10299 1643 10699
rect 2033 10299 2038 10699
rect 1638 10294 2038 10299
rect 480 840 31720 880
rect 480 520 520 840
rect 840 520 31360 840
rect 31680 520 31720 840
rect 480 480 31720 520
rect 0 360 32200 400
rect 0 40 40 360
rect 360 40 31840 360
rect 32160 40 32200 360
rect 0 0 32200 40
<< via3 >>
rect 28832 21842 28896 21906
rect 31897 21728 32073 21733
rect 31897 21552 31902 21728
rect 31902 21552 32068 21728
rect 32068 21552 32073 21728
rect 31897 21547 32073 21552
rect 31381 20788 31557 20793
rect 31381 20612 31386 20788
rect 31386 20612 31552 20788
rect 31552 20612 31557 20788
rect 31381 20607 31557 20612
rect 31802 13534 32200 13934
rect 31323 12823 31721 13223
rect 0 11036 398 11436
rect 479 10299 877 10699
rect 520 520 840 840
rect 31360 520 31680 840
rect 40 40 360 360
rect 31840 40 32160 360
<< metal4 >>
rect 0 11437 400 22304
rect -1 11436 400 11437
rect -1 11036 0 11436
rect 398 11036 400 11436
rect -1 11035 400 11036
rect 0 360 400 11035
rect 480 10700 880 22304
rect 6134 22104 6194 22304
rect 6686 22104 6746 22304
rect 7238 22104 7298 22304
rect 7790 19852 7850 22304
rect 8342 22104 8402 22304
rect 8894 22104 8954 22304
rect 9446 22104 9506 22304
rect 9998 22104 10058 22304
rect 10550 22104 10610 22304
rect 11102 22104 11162 22304
rect 11654 22104 11714 22304
rect 12206 22104 12266 22304
rect 12758 22104 12818 22304
rect 13310 22104 13370 22304
rect 13862 22104 13922 22304
rect 14414 22104 14474 22304
rect 14966 22104 15026 22304
rect 15518 22104 15578 22304
rect 16070 22104 16130 22304
rect 16622 19840 16682 22304
rect 17174 22046 17234 22304
rect 17726 22046 17786 22304
rect 18278 22046 18338 22304
rect 18830 22046 18890 22304
rect 19382 22046 19442 22304
rect 19934 22046 19994 22304
rect 20486 22046 20546 22304
rect 21038 22104 21098 22304
rect 21590 22104 21650 22304
rect 22142 22104 22202 22304
rect 22694 22104 22754 22304
rect 23246 22104 23306 22304
rect 23798 22104 23858 22304
rect 24350 22104 24410 22304
rect 24902 22104 24962 22304
rect 25454 22034 25514 22304
rect 25454 21920 25514 21974
rect 26006 22038 26066 22304
rect 26006 21920 26066 21978
rect 26558 22024 26618 22304
rect 26558 21920 26618 21964
rect 27110 22032 27170 22304
rect 27110 21920 27170 21972
rect 27662 22038 27722 22304
rect 27662 21920 27722 21978
rect 28214 22034 28274 22304
rect 28214 21920 28274 21974
rect 28766 22036 28826 22304
rect 28766 21920 28826 21976
rect 29318 22032 29378 22304
rect 29318 21920 29378 21972
rect 25382 21906 29378 21920
rect 25382 21848 28832 21906
rect 28831 21842 28832 21848
rect 28896 21870 29378 21906
rect 28896 21848 29372 21870
rect 28896 21842 28897 21848
rect 28831 21841 28897 21842
rect 31320 20793 31720 22304
rect 31320 20607 31381 20793
rect 31557 20607 31720 20793
rect 478 10699 880 10700
rect 478 10299 479 10699
rect 877 10299 880 10699
rect 478 10298 880 10299
rect 0 40 40 360
rect 360 40 400 360
rect 0 0 400 40
rect 480 840 880 10298
rect 480 520 520 840
rect 840 520 880 840
rect 480 0 880 520
rect 31320 13224 31720 20607
rect 31800 21733 32200 22304
rect 31800 21547 31897 21733
rect 32073 21547 32200 21733
rect 31800 13935 32200 21547
rect 31800 13934 32201 13935
rect 31800 13534 31802 13934
rect 32200 13534 32201 13934
rect 31800 13533 32201 13534
rect 31320 13223 31722 13224
rect 31320 12823 31323 13223
rect 31721 12823 31722 13223
rect 31320 12822 31722 12823
rect 31320 840 31720 12822
rect 31320 520 31360 840
rect 31680 520 31720 840
rect 31320 0 31720 520
rect 31800 360 32200 13533
rect 31800 40 31840 360
rect 32160 40 32200 360
rect 31800 0 32200 40
<< rmetal4 >>
rect 25454 21974 25514 22034
rect 26006 21978 26066 22038
rect 26558 21964 26618 22024
rect 27110 21972 27170 22032
rect 27662 21978 27722 22038
rect 28214 21974 28274 22034
rect 28766 21976 28826 22036
rect 29318 21972 29378 22032
use JNWTR_TAPCELLB_CV  JNWTR_TAPCELLB_CV_0 JNW_TR_SKY130A
timestamp 1769070524
transform 1 0 27886 0 1 20846
box -150 -120 2130 440
use JNWTR_TIEL_CV  JNWTR_TIEL_CV_0 JNW_TR_SKY130A
timestamp 1769070524
transform 1 0 27886 0 1 21166
box -150 -120 2130 440
use LELO_GR02  LELO_GR02_0
timestamp 1769081024
transform 1 0 1100 0 1 1200
box 0 0 30000 19000
<< labels >>
flabel metal4 s 6686 22104 6746 22304 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 6134 22104 6194 22304 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 7238 22104 7298 22304 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 7790 22104 7850 22304 0 FreeSans 480 90 0 0 ui_in[0]
port 3 nsew signal input
flabel metal4 s 8342 22104 8402 22304 0 FreeSans 480 90 0 0 ui_in[1]
port 4 nsew signal input
flabel metal4 s 8894 22104 8954 22304 0 FreeSans 480 90 0 0 ui_in[2]
port 5 nsew signal input
flabel metal4 s 9446 22104 9506 22304 0 FreeSans 480 90 0 0 ui_in[3]
port 6 nsew signal input
flabel metal4 s 9998 22104 10058 22304 0 FreeSans 480 90 0 0 ui_in[4]
port 7 nsew signal input
flabel metal4 s 10550 22104 10610 22304 0 FreeSans 480 90 0 0 ui_in[5]
port 8 nsew signal input
flabel metal4 s 11102 22104 11162 22304 0 FreeSans 480 90 0 0 ui_in[6]
port 9 nsew signal input
flabel metal4 s 11654 22104 11714 22304 0 FreeSans 480 90 0 0 ui_in[7]
port 10 nsew signal input
flabel metal4 s 12206 22104 12266 22304 0 FreeSans 480 90 0 0 uio_in[0]
port 11 nsew signal input
flabel metal4 s 12758 22104 12818 22304 0 FreeSans 480 90 0 0 uio_in[1]
port 12 nsew signal input
flabel metal4 s 13310 22104 13370 22304 0 FreeSans 480 90 0 0 uio_in[2]
port 13 nsew signal input
flabel metal4 s 13862 22104 13922 22304 0 FreeSans 480 90 0 0 uio_in[3]
port 14 nsew signal input
flabel metal4 s 14414 22104 14474 22304 0 FreeSans 480 90 0 0 uio_in[4]
port 15 nsew signal input
flabel metal4 s 14966 22104 15026 22304 0 FreeSans 480 90 0 0 uio_in[5]
port 16 nsew signal input
flabel metal4 s 15518 22104 15578 22304 0 FreeSans 480 90 0 0 uio_in[6]
port 17 nsew signal input
flabel metal4 s 16070 22104 16130 22304 0 FreeSans 480 90 0 0 uio_in[7]
port 18 nsew signal input
flabel metal4 s 25454 22104 25514 22304 0 FreeSans 480 90 0 0 uio_oe[0]
port 19 nsew signal output
flabel metal4 s 26006 22104 26066 22304 0 FreeSans 480 90 0 0 uio_oe[1]
port 20 nsew signal output
flabel metal4 s 26558 22104 26618 22304 0 FreeSans 480 90 0 0 uio_oe[2]
port 21 nsew signal output
flabel metal4 s 27110 22104 27170 22304 0 FreeSans 480 90 0 0 uio_oe[3]
port 22 nsew signal output
flabel metal4 s 27662 22104 27722 22304 0 FreeSans 480 90 0 0 uio_oe[4]
port 23 nsew signal output
flabel metal4 s 28214 22104 28274 22304 0 FreeSans 480 90 0 0 uio_oe[5]
port 24 nsew signal output
flabel metal4 s 28766 22104 28826 22304 0 FreeSans 480 90 0 0 uio_oe[6]
port 25 nsew signal output
flabel metal4 s 21038 22104 21098 22304 0 FreeSans 480 90 0 0 uio_out[0]
port 27 nsew signal output
flabel metal4 s 21590 22104 21650 22304 0 FreeSans 480 90 0 0 uio_out[1]
port 28 nsew signal output
flabel metal4 s 22142 22104 22202 22304 0 FreeSans 480 90 0 0 uio_out[2]
port 29 nsew signal output
flabel metal4 s 22694 22104 22754 22304 0 FreeSans 480 90 0 0 uio_out[3]
port 30 nsew signal output
flabel metal4 s 23246 22104 23306 22304 0 FreeSans 480 90 0 0 uio_out[4]
port 31 nsew signal output
flabel metal4 s 23798 22104 23858 22304 0 FreeSans 480 90 0 0 uio_out[5]
port 32 nsew signal output
flabel metal4 s 24350 22104 24410 22304 0 FreeSans 480 90 0 0 uio_out[6]
port 33 nsew signal output
flabel metal4 s 24902 22104 24962 22304 0 FreeSans 480 90 0 0 uio_out[7]
port 34 nsew signal output
flabel metal4 s 16622 22104 16682 22304 0 FreeSans 480 90 0 0 uo_out[0]
port 35 nsew signal output
flabel metal4 s 17174 22104 17234 22304 0 FreeSans 480 90 0 0 uo_out[1]
port 36 nsew signal output
flabel metal4 s 17726 22104 17786 22304 0 FreeSans 480 90 0 0 uo_out[2]
port 37 nsew signal output
flabel metal4 s 18278 22104 18338 22304 0 FreeSans 480 90 0 0 uo_out[3]
port 38 nsew signal output
flabel metal4 s 18830 22104 18890 22304 0 FreeSans 480 90 0 0 uo_out[4]
port 39 nsew signal output
flabel metal4 s 19382 22104 19442 22304 0 FreeSans 480 90 0 0 uo_out[5]
port 40 nsew signal output
flabel metal4 s 19934 22104 19994 22304 0 FreeSans 480 90 0 0 uo_out[6]
port 41 nsew signal output
flabel metal4 s 20486 22104 20546 22304 0 FreeSans 480 90 0 0 uo_out[7]
port 42 nsew signal output
flabel metal4 480 0 880 22304 1 FreeSans 800 0 0 0 VGND
port 44 nsew ground bidirectional
flabel metal4 0 0 400 22304 1 FreeSans 800 0 0 0 VDPWR
port 43 nsew power bidirectional
flabel metal4 s 29318 22104 29378 22304 0 FreeSans 480 90 0 0 uio_oe[7]
port 26 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 32200 22304
<< end >>
