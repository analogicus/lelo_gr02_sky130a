*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/BANDGAP_OPAMP_lpe.spi
#else
.include ../../../work/xsch/BANDGAP_OPAMP.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p
.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS    VSS       0    dc 0
VDD    VDD_1V8   VSS  pwl 0 0 5n {AVDD}
VPWR  PWRUP_1V8  VSS  dc 0
V_POS  VIN_N     VSS  dc 0.5 ac 0.5 sin(0 0.5 100MEG)  
V_NEG  VIN_P     VSS  dc 0.5
*---------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save all

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 1u 0


tran 1n 300n 1p
write
quit


.endc

.end
