** sch_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/BANDGAP_OPAMP/BANDGAP_OPAMP.sch
**.subckt BANDGAP_OPAMP VDD_1V8 PWRUP_1V8 VOUT VIN_N VIN_P VSS
*.ipin VDD_1V8
*.ipin VSS
*.ipin PWRUP_1V8
*.ipin VIN_P
*.ipin VIN_N
*.opin VOUT
x8 SUPPLY PWRUP_1V8 VDD_1V8 VDD_1V8 JNWATR_PCH_12C1F2
R1 SUPPLY V_IB 100k m=1
x5<5> PMOS_GATE VIN_P TAIL VSS JNWATR_NCH_4C1F2
x5<4> PMOS_GATE VIN_P TAIL VSS JNWATR_NCH_4C1F2
x5<3> PMOS_GATE VIN_P TAIL VSS JNWATR_NCH_4C1F2
x5<2> PMOS_GATE VIN_P TAIL VSS JNWATR_NCH_4C1F2
x5<1> PMOS_GATE VIN_P TAIL VSS JNWATR_NCH_4C1F2
x5<0> PMOS_GATE VIN_P TAIL VSS JNWATR_NCH_4C1F2
x3<5> net1 VIN_N TAIL VSS JNWATR_NCH_4C1F2
x3<4> net1 VIN_N TAIL VSS JNWATR_NCH_4C1F2
x3<3> net1 VIN_N TAIL VSS JNWATR_NCH_4C1F2
x3<2> net1 VIN_N TAIL VSS JNWATR_NCH_4C1F2
x3<1> net1 VIN_N TAIL VSS JNWATR_NCH_4C1F2
x3<0> net1 VIN_N TAIL VSS JNWATR_NCH_4C1F2
x4 V_IB V_IB VSS VSS JNWATR_NCH_4C1F2
x6 TAIL V_IB VSS VSS JNWATR_NCH_4C1F2
x7 net1 PMOS_GATE SUPPLY VDD_1V8 JNWATR_PCH_4C1F2
x1 PMOS_GATE PMOS_GATE SUPPLY VDD_1V8 JNWATR_PCH_4C1F2
x2 VOUT net1 SUPPLY VDD_1V8 JNWATR_PCH_4C1F2
x3 VOUT V_IB VSS VSS JNWATR_NCH_4C1F2
**.ends

* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_PCH_12C1F2.sym # of pins=4
** sym_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_12C1F2.sym
** sch_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_12C1F2.sch
.subckt JNWATR_PCH_12C1F2 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.22 W=8.32 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_NCH_4C1F2.sym # of pins=4
** sym_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_4C1F2.sym
** sch_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_4C1F2.sch
.subckt JNWATR_NCH_4C1F2 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.22 W=3.2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_PCH_4C1F2.sym # of pins=4
** sym_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C1F2.sym
** sch_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C1F2.sch
.subckt JNWATR_PCH_4C1F2 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.22 W=3.2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
