** sch_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/LELO_GR02_SKY130A/TB_LELOGR02_BANDGAP_OPAMP.sch
**.subckt TB_LELOGR02_BANDGAP_OPAMP
V1 TB_VIP 0 sin(0.8 0.5m 10k)
V2 TB_VIN 0 sin(0.8 -0.5m 10k)
x5 TB_VOUT 0 JNWTR_CAPX1
V3 TB_VDD 0 1.8
x1 TB_VDD 0 TB_VOUT TB_VIN TB_VIP 0 OPAMP2
**** begin user architecture code


.param mc_mm_switch=0
.param mc_pr_switch=0

.lib ../../../tech/ngspice/temperature.spi Tl
.lib ../../../tech/ngspice/corners.spi Kss
.lib ../../../tech/ngspice/supply.spi Vl
.include ../../../../cpdk/ngspice/ideal_circuits.spi

.option SEED=1
.option savevoltages
.option gmin=1e-12
.control


optran 0 0 0 10n 1u 0
op
write TB_OPAMP2_op.raw

*tran 1u 200u
*write TB_OPAMP2_tran.raw



exit
.endc



**** end user architecture code
**.ends

* expanding   symbol:  JNW_TR_SKY130A/JNWTR_CAPX1.sym # of pins=2
** sym_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_CAPX1.sym
** sch_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_CAPX1.sch
.subckt JNWTR_CAPX1 A B
*.iopin A
*.iopin B
XC1 B A sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
.ends


* expanding   symbol:  OPAMP2.sym # of pins=6
** sym_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/OPAMP2.sym
** sch_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/OPAMP2.sch
.subckt OPAMP2 VDD_1V8 PWRUP_1V8 VOUT VIN_N VIN_P VSS
*.ipin VDD_1V8
*.ipin VSS
*.ipin PWRUP_1V8
*.ipin VIN_P
*.opin VOUT
*.ipin VIN_N
x8 SUPPLY PWRUP_1V8 VDD_1V8 VDD_1V8 JNWATR_PCH_2C1F2
x2 V_IB net2 VSS JNWTR_RPPO16
x7 V_IB V_IB VSS VSS JNWATR_NCH_4C5F0
x3 TAIL V_IB VSS VSS JNWATR_NCH_4C5F0
x4<3> VOUT V_IB VSS VSS JNWATR_NCH_4C5F0
x4<2> VOUT V_IB VSS VSS JNWATR_NCH_4C5F0
x4<1> VOUT V_IB VSS VSS JNWATR_NCH_4C5F0
x4<0> VOUT V_IB VSS VSS JNWATR_NCH_4C5F0
x10<4> net1 VIN_P TAIL VSS LELOATR_LVT_NCH_4C5F0
x10<3> net1 VIN_P TAIL VSS LELOATR_LVT_NCH_4C5F0
x10<2> net1 VIN_P TAIL VSS LELOATR_LVT_NCH_4C5F0
x10<1> net1 VIN_P TAIL VSS LELOATR_LVT_NCH_4C5F0
x10<0> net1 VIN_P TAIL VSS LELOATR_LVT_NCH_4C5F0
x1<4> PMOS_GATE VIN_N TAIL VSS LELOATR_LVT_NCH_4C5F0
x1<3> PMOS_GATE VIN_N TAIL VSS LELOATR_LVT_NCH_4C5F0
x1<2> PMOS_GATE VIN_N TAIL VSS LELOATR_LVT_NCH_4C5F0
x1<1> PMOS_GATE VIN_N TAIL VSS LELOATR_LVT_NCH_4C5F0
x1<0> PMOS_GATE VIN_N TAIL VSS LELOATR_LVT_NCH_4C5F0
x6 net1 PMOS_GATE SUPPLY VDD_1V8 JNWATR_PCH_4C5F0
x11 PMOS_GATE PMOS_GATE SUPPLY VDD_1V8 JNWATR_PCH_4C5F0
x2<5> net1 VOUT JNWTR_CAPX4
x2<4> net1 VOUT JNWTR_CAPX4
x2<3> net1 VOUT JNWTR_CAPX4
x2<2> net1 VOUT JNWTR_CAPX4
x2<1> net1 VOUT JNWTR_CAPX4
x2<0> net1 VOUT JNWTR_CAPX4
x3<3> VOUT net1 SUPPLY VDD_1V8 LELOATR_LVT_PCH_4C5F0
x3<2> VOUT net1 SUPPLY VDD_1V8 LELOATR_LVT_PCH_4C5F0
x3<1> VOUT net1 SUPPLY VDD_1V8 LELOATR_LVT_PCH_4C5F0
x3<0> VOUT net1 SUPPLY VDD_1V8 LELOATR_LVT_PCH_4C5F0
x9 net2 SUPPLY VSS JNWTR_RPPO16
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_PCH_2C1F2.sym # of pins=4
** sym_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_2C1F2.sym
** sch_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_2C1F2.sch
.subckt JNWATR_PCH_2C1F2 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.22 W=1.92 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RPPO16.sym # of pins=3
** sym_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO16.sym
** sch_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO16.sch
.subckt JNWTR_RPPO16 N P B
*.iopin P
*.iopin N
*.iopin B
XXA1 N P B JNWTR_RES16
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sym # of pins=4
** sym_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sym
** sch_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sch
.subckt JNWATR_NCH_4C5F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.94 W=3.2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  LELO_ATR_SKY130A/LELOATR_LVT_NCH_4C5F0.sym # of pins=4
** sym_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/LELO_ATR_SKY130A/LELOATR_LVT_NCH_4C5F0.sym
** sch_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/LELO_ATR_SKY130A/LELOATR_LVT_NCH_4C5F0.sch
.subckt LELOATR_LVT_NCH_4C5F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8_lvt L=0.94 W=3.2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_PCH_4C5F0.sym # of pins=4
** sym_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C5F0.sym
** sch_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C5F0.sch
.subckt JNWATR_PCH_4C5F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.94 W=3.2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_CAPX4.sym # of pins=2
** sym_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_CAPX4.sym
** sch_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_CAPX4.sch
.subckt JNWTR_CAPX4 A B
*.iopin A
*.iopin B
XXA1 A B JNWTR_CAPX1
XXA2 A B JNWTR_CAPX1
XXB1 A B JNWTR_CAPX1
XXB2 A B JNWTR_CAPX1
.ends


* expanding   symbol:  LELO_ATR_SKY130A/LELOATR_LVT_PCH_4C5F0.sym # of pins=4
** sym_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/LELO_ATR_SKY130A/LELOATR_LVT_PCH_4C5F0.sym
** sch_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/LELO_ATR_SKY130A/LELOATR_LVT_PCH_4C5F0.sch
.subckt LELOATR_LVT_PCH_4C5F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8_lvt L=0.94 W=3.2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RES16.sym # of pins=3
** sym_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RES16.sym
** sch_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_RES16.sch
.subckt JNWTR_RES16 N P B
*.iopin N
*.iopin P
*.iopin B
XR1_0 INT_0 N B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_1 INT_1 INT_0 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_2 INT_2 INT_1 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_3 INT_3 INT_2 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_4 INT_4 INT_3 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_5 INT_5 INT_4 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_6 INT_6 INT_5 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_7 INT_7 INT_6 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_8 INT_8 INT_7 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_9 INT_9 INT_8 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_10 INT_10 INT_9 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_11 INT_11 INT_10 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_12 INT_12 INT_11 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_13 INT_13 INT_12 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_14 INT_14 INT_13 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_15 P INT_14 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
.ends

.end
