** sch_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/LELO_GR02_SKY130A/TB_OPAMP.sch
**.subckt TB_OPAMP
V1 net1 0 1.8
.save i(v1)
V2 VIN_N 0 sin(0.7 50m 10k)
V3 VIN_P 0 0.7
x5 VOUT 0 JNWTR_CAPX1
x1 net1 0 VOUT VIN_N VIN_P 0 BANDGAP_OPAMP
**** begin user architecture code


.param mc_mm_switch=0
.param mc_pr_switch=0

.lib /home/ivera/pro/aicex/ip/tech_sky130A/ngspice/temperature.spi Tl
.lib /home/ivera/pro/aicex/ip/tech_sky130A/ngspice/corners.spi Kss
.lib /home/ivera/pro/aicex/ip/tech_sky130A/ngspice/supply.spi Vl
.include /home/ivera/pro/aicex/ip/cpdk/ngspice/ideal_circuits.spi

.option SEED=1
.option savecurrents
.save all
.control

optran 0 0 0 10n 1u 0


tran 100n 200u
write TB_graph.raw

*exit
.endc



**** end user architecture code
**.ends

* expanding   symbol:  JNW_TR_SKY130A/JNWTR_CAPX1.sym # of pins=2
** sym_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_CAPX1.sym
** sch_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_TR_SKY130A/JNWTR_CAPX1.sch
.subckt JNWTR_CAPX1 A B
*.iopin A
*.iopin B
XC1 B A sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
.ends


* expanding   symbol:  BANDGAP_OPAMP/BANDGAP_OPAMP.sym # of pins=6
** sym_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/BANDGAP_OPAMP/BANDGAP_OPAMP.sym
** sch_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/BANDGAP_OPAMP/BANDGAP_OPAMP.sch
.subckt BANDGAP_OPAMP VDD_1V8 PWRUP_1V8 VOUT VIN_N VIN_P VSS
*.ipin VDD_1V8
*.ipin VSS
*.ipin PWRUP_1V8
*.ipin VIN_P
*.ipin VIN_N
*.opin VOUT
x3 net1 VIN_P net2 VSS JNWATR_NCH_4C5F0
x4 VOUT VIN_N net2 VSS JNWATR_NCH_4C5F0
x1 VOUT net1 net4 net4 JNWATR_PCH_4C5F0
x2 net1 net1 net4 net4 JNWATR_PCH_4C5F0
x6 net5 net3 VSS VSS JNWATR_NCH_4C5F0
x7 net2 net3 VSS VSS JNWATR_NCH_4C5F0
x8 net4 PWRUP_1V8 VDD_1V8 VDD_1V8 JNWATR_PCH_12C1F2
R1 net5 net4 sky130_fd_pr__res_generic_m4 W=1 L=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sym # of pins=4
** sym_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sym
** sch_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sch
.subckt JNWATR_NCH_4C5F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.94 W=3.2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_PCH_4C5F0.sym # of pins=4
** sym_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C5F0.sym
** sch_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C5F0.sch
.subckt JNWATR_PCH_4C5F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.94 W=3.2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_PCH_12C1F2.sym # of pins=4
** sym_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_12C1F2.sym
** sch_path: /home/ivera/pro/aicex/ip/lelo_gr02_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_12C1F2.sch
.subckt JNWATR_PCH_12C1F2 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.22 W=8.32 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
