*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/BANDGAP_OPAMP_lpe.spi
#else
.include ../../../work/xsch/BANDGAP_OPAMP.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p
.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS    VSS       0    dc 0
VDD    VDD_1V8   VSS  dc {AVDD}
VPWR   PWRUP_1V8 VSS  dc pwl(0 {AVDD}, 50n {AVDD}, 50.1n 0)
V_POS  VIP       VSS  dc sin(0.5 0.5m 10k)  
V_NEG  VIN       VSS  dc 0.5
*---------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save all

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 1u 0


tran 1u 100m 1p
write
quit


.endc

.end
